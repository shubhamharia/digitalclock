----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 15.03.2021 20:33:04
-- Design Name: 
-- Module Name: clockdivide_tb - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity multiplexer_tb is
--  Port ( );
end multiplexer_tb;

architecture Behavioral of multiplexer_tb is
component multiplexer is 
  Port ( clockin : in STD_LOGIC;
           sel : out STD_LOGIC_VECTOR (1 downto 0));
end component;
--input
signal clockin:STD_LOGIC:='0';
--OUTPUR
signal sel: STD_LOGIC_VECTOR (1 downto 0);
constant clk_period : time :=100 ns;

begin
utt:multiplexer  port map(
clockin=> clockin,
sel=>sel);
timer:process
begin
clockin<='1';
wait for clk_period/2;
clockin<='0';
wait for clk_period/2;
end process;
end Behavioral;

